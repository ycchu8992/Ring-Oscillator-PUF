`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:
// Design Name: 
// Module Name: scrambler
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: scrambler_lfsr builds on top of the existing LFSR module and adds
//             an element on nonlinearity to it making it harder to predict.
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module scrambler(input_challenge, clk, rst, output_challenge);
input [7:0] input_challenge;
input clk, rst;
output reg [7:0] output_challenge;

***************
**Your Coding**
***************

endmodule
