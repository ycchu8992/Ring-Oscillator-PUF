`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 
// Design Name: 
// Module Name: MUX_8to1
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: The MUX_8to1 is a multiplexer that selects between 8 inputs
//               and passes through only one. It follows that the select line
//               is a 4-bit bus.
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module MUX_8to1(a,b,c,d,e,f,g,h,sel,mux_out);
input a,b,c,d,e,f,g,h;
input [3:0] sel;	//from the output of scrambler
output reg mux_out;

***************
**Your Coding**
***************

endmodule
